`timescale 1ns / 1ps

module wrapper_tb;

    reg         clk;
    reg         reset;
    reg         reset2;
    reg [11:0]   address;
    reg [63:0]  writedata;
    reg         write;
    reg         read;
    reg [7:0] byteenable;
    wire [63:0] readdata;
    wire        waitrequest;

    avalonsuxx dut_inst(clk, reset, address, writedata, write, read, byteenable, readdata, waitrequest);

    always begin
        #5 clk <= ~clk;
    end

    initial begin
        clk = 1; reset = 1; reset2 = 1;
        #20 reset = 0; reset2 = 0;   
        #10 address =  0 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  3 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  4 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  5 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  6 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  7 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  8 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  9 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  10 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  11 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  12 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  13 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  14 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  15 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  16 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  17 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  18 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  19 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  20 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  21 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  22 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  23 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  24 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  25 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  26 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  27 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  28 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  29 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  30 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  31 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  32 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  33 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  34 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  35 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  36 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  37 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  38 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  39 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  40 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  41 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  42 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  43 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  44 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  45 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  46 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  47 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  48 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  49 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  50 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  51 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  52 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  53 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  54 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  55 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  56 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  57 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  58 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  59 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  60 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  61 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  62 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  63 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  64 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  65 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  66 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  67 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  68 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  69 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  70 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  71 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  72 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  73 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  74 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  75 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  76 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  77 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  78 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  79 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  80 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  81 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  82 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  83 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  84 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  85 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  86 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  87 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  88 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  89 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  90 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  91 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  92 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  93 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  94 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  95 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  96 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  97 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  98 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  99 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  100 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  101 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  102 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  103 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  104 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  105 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  106 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  107 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  108 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  109 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  110 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  111 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  112 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  113 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  114 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  115 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  116 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  117 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  118 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  119 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  120 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  121 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  122 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  123 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  124 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  125 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  126 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  127 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  128 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  129 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  130 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  131 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  132 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  133 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  134 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  135 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  136 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  137 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  138 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  139 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  140 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  141 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  142 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  143 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  144 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  145 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  146 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  147 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  148 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  149 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  150 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  151 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  152 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  153 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  154 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  155 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  156 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  157 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  158 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  159 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  160 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  161 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  162 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  163 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  164 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  165 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  166 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  167 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  168 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  169 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  170 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  171 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  172 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  173 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  174 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  175 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  176 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  177 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  178 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  179 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  180 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  181 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  182 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  183 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  184 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  185 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  186 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  187 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  188 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  189 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  190 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  191 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  192 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  193 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  194 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  195 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  196 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  197 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  198 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  199 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  200 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  201 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  202 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  203 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  204 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  205 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  206 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  207 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  208 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  209 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  210 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  211 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  212 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  213 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  214 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  215 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  216 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  217 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  218 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  219 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  220 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  221 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  222 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  223 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  224 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  225 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  226 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  227 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  228 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  229 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  230 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  231 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  232 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  233 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  234 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  235 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  236 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  237 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  238 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  239 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  240 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  241 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  242 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  243 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  244 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  245 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  246 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  247 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  248 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  249 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  250 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  251 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  252 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  253 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  254 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  255 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  256 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  257 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  258 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  259 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  260 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  261 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  262 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  263 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  264 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  265 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  266 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  267 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  268 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  269 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  270 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  271 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  272 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  273 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  274 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  275 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  276 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  277 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  278 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  279 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  280 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  281 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  282 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  283 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  284 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  285 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  286 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  287 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  288 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  289 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  290 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  291 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  292 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  293 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  294 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  295 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  296 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  297 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  298 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  299 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  300 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  301 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  302 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  303 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  304 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  305 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  306 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  307 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  308 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  309 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  310 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  311 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  312 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  313 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  314 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  315 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  316 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  317 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  318 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  319 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  320 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  321 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  322 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  323 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  324 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  325 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  326 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  327 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  328 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  329 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  330 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  331 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  332 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  333 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  334 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  335 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  336 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  337 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  338 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  339 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  340 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  341 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  342 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  343 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  344 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  345 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  346 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  347 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  348 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  349 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  350 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  351 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  352 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  353 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  354 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  355 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  356 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  357 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  358 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  359 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  360 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  361 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  362 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  363 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  364 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  365 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  366 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  367 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  368 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  369 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  370 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  371 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  372 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  373 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  374 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  375 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  376 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  377 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  378 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  379 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  380 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  381 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  382 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  383 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  384 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  385 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  386 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  387 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  388 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  389 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  390 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  391 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  392 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  393 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  394 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  395 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  396 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  397 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  398 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  399 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  400 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  401 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  402 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  403 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  404 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  405 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  406 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  407 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  408 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  409 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  410 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  411 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  412 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  413 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  414 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  415 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  416 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  417 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  418 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  419 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  420 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  421 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  422 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  423 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  424 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  425 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  426 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  427 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  428 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  429 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  430 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  431 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  432 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  433 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  434 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  435 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  436 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  437 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  438 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  439 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  440 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  441 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  442 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  443 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  444 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  445 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  446 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  447 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  448 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  449 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  450 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  451 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  452 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  453 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  454 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  455 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  456 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  457 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  458 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  459 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  460 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  461 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  462 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  463 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  464 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  465 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  466 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  467 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  468 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  469 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  470 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  471 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  472 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  473 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  474 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  475 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  476 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  477 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  478 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  479 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  480 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  481 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  482 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  483 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  484 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  485 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  486 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  487 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  488 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  489 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  490 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  491 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  492 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  493 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  494 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  495 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  496 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  497 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  498 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  499 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  500 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  501 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  502 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  503 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  504 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  505 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  506 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  507 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  508 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  509 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  510 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  511 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  512 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  513 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  514 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  515 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  516 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  517 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  518 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  519 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  520 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  521 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  522 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  523 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  524 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  525 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  526 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  527 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  528 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  529 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  530 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  531 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  532 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  533 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  534 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  535 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  536 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  537 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  538 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  539 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  540 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  541 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  542 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  543 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  544 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  545 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  546 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  547 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  548 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  549 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  550 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  551 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  552 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  553 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  554 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  555 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  556 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  557 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  558 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  559 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  560 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  561 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  562 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  563 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  564 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  565 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  566 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  567 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  568 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  569 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  570 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  571 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  572 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  573 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  574 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  575 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  576 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  577 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  578 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  579 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  580 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  581 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  582 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  583 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  584 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  585 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  586 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  587 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  588 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  589 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  590 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  591 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  592 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  593 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  594 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  595 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  596 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  597 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  598 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  599 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  600 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  601 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  602 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  603 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  604 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  605 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  606 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  607 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  608 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  609 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  610 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  611 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  612 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  613 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  614 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  615 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  616 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  617 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  618 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  619 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  620 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  621 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  622 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  623 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  624 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  625 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  626 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  627 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  628 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  629 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  630 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  631 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  632 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  633 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  634 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  635 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  636 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  637 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  638 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  639 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  640 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  641 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  642 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  643 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  644 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  645 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  646 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  647 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  648 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  649 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  650 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  651 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  652 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  653 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  654 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  655 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  656 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  657 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  658 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  659 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  660 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  661 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  662 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  663 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  664 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  665 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  666 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  667 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  668 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  669 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  670 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  671 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  672 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  673 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  674 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  675 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  676 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  677 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  678 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  679 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  680 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  681 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  682 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  683 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  684 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  685 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  686 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  687 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  688 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  689 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  690 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  691 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  692 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  693 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  694 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  695 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  696 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  697 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  698 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  699 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  700 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  701 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  702 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  703 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  704 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  705 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  706 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  707 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  708 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  709 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  710 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  711 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  712 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  713 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  714 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  715 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  716 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  717 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  718 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  719 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  720 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  721 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  722 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  723 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  724 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  725 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  726 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  727 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  728 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  729 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  730 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  731 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  732 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  733 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  734 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  735 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  736 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  737 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  738 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  739 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  740 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  741 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  742 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  743 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  744 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  745 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  746 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  747 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  748 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  749 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  750 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  751 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  752 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  753 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  754 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  755 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  756 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  757 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  758 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  759 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  760 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  761 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  762 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  763 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  764 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  765 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  766 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  767 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  768 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  769 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  770 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  771 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  772 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  773 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  774 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  775 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  776 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  777 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  778 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  779 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  780 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  781 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  782 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  783 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  784 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  785 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  786 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  787 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  788 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  789 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  790 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  791 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  792 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  793 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  794 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  795 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  796 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  797 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  798 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  799 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  800 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  801 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  802 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  803 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  804 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  805 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  806 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  807 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  808 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  809 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  810 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  811 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  812 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  813 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  814 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  815 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  816 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  817 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  818 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  819 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  820 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  821 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  822 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  823 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  824 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  825 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  826 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  827 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  828 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  829 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  830 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  831 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  832 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  833 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  834 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  835 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  836 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  837 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  838 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  839 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  840 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  841 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  842 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  843 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  844 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  845 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  846 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  847 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  848 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  849 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  850 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  851 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  852 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  853 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  854 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  855 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  856 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  857 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  858 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  859 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  860 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  861 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  862 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  863 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  864 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  865 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  866 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  867 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  868 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  869 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  870 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  871 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  872 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  873 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  874 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  875 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  876 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  877 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  878 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  879 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  880 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  881 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  882 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  883 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  884 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  885 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  886 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  887 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  888 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  889 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  890 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  891 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  892 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  893 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  894 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  895 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  896 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  897 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  898 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  899 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  900 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  901 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  902 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  903 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  904 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  905 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  906 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  907 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  908 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  909 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  910 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  911 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  912 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  913 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  914 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  915 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  916 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  917 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  918 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  919 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  920 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  921 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  922 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  923 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  924 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  925 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  926 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  927 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  928 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  929 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  930 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  931 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  932 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  933 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  934 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  935 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  936 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  937 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  938 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  939 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  940 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  941 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  942 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  943 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  944 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  945 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  946 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  947 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  948 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  949 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  950 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  951 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  952 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  953 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  954 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  955 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  956 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  957 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  958 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  959 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  960 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  961 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  962 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  963 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  964 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  965 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  966 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  967 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  968 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  969 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  970 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  971 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  972 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  973 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  974 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  975 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  976 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  977 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  978 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  979 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  980 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  981 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  982 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  983 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  984 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  985 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  986 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  987 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  988 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  989 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  990 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  991 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  992 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  993 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  994 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  995 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  996 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  997 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  998 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  999 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1000 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1001 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1002 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1003 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1004 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1005 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1006 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1007 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1008 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1009 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1010 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1011 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1012 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1013 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1014 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1015 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1016 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1017 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1018 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1019 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1020 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1021 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1022 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1023 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1024 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1025 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1026 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1027 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1028 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1029 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1030 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1031 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1032 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1033 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1034 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1035 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1036 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1037 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1038 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1039 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1040 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1041 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1042 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1043 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1044 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1045 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1046 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1047 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1048 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1049 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1050 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1051 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1052 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1053 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1054 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1055 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1056 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1057 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1058 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1059 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1060 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1061 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1062 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1063 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1064 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1065 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1066 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1067 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1068 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1069 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1070 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1071 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1072 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1073 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1074 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1075 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1076 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1077 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1078 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1079 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1080 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1081 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1082 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1083 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1084 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1085 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1086 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1087 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1088 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1089 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1090 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1091 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1092 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1093 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1094 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1095 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1096 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1097 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1098 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1099 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1100 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1101 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1102 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1103 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1104 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1105 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1106 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1107 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1108 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1109 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1110 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1111 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1112 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1113 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1114 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1115 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1116 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1117 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1118 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1119 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1120 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1121 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1122 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1123 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1124 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1125 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1126 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1127 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1128 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1129 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1130 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1131 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1132 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1133 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1134 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1135 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1136 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1137 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1138 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1139 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1140 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1141 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1142 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1143 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1144 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1145 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1146 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1147 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1148 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1149 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1150 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1151 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1152 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1153 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1154 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1155 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1156 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1157 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1158 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1159 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1160 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1161 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1162 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1163 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1164 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1165 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1166 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1167 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1168 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1169 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1170 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1171 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1172 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1173 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1174 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1175 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1176 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1177 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1178 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1179 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1180 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1181 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1182 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1183 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1184 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1185 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1186 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1187 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1188 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1189 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1190 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1191 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1192 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1193 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1194 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1195 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1196 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1197 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1198 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1199 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1200 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1201 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1202 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1203 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1204 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1205 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1206 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1207 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1208 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1209 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1210 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1211 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1212 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1213 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1214 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1215 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1216 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1217 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1218 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1219 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1220 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1221 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1222 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1223 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1224 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1225 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1226 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1227 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1228 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1229 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1230 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1231 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1232 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1233 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1234 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1235 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1236 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1237 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1238 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1239 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1240 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1241 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1242 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1243 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1244 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1245 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1246 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1247 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1248 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1249 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1250 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1251 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1252 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1253 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1254 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1255 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1256 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1257 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1258 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1259 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1260 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1261 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1262 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1263 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1264 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1265 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1266 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1267 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1268 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1269 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1270 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1271 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1272 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1273 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1274 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1275 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1276 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1277 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1278 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1279 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1280 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1281 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1282 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1283 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1284 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1285 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1286 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1287 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1288 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1289 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1290 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1291 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1292 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1293 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1294 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1295 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1296 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1297 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1298 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1299 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1300 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1301 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1302 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1303 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1304 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1305 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1306 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1307 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1308 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1309 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1310 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1311 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1312 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1313 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1314 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1315 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1316 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1317 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1318 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1319 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1320 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1321 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1322 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1323 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1324 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1325 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1326 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1327 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1328 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1329 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1330 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1331 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1332 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1333 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1334 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1335 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1336 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1337 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1338 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1339 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1340 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1341 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1342 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1343 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1344 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1345 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1346 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1347 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1348 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1349 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1350 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1351 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1352 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1353 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1354 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1355 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1356 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1357 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1358 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1359 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1360 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1361 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1362 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1363 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1364 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1365 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1366 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1367 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1368 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1369 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1370 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1371 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1372 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1373 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1374 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1375 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1376 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1377 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1378 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1379 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1380 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1381 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1382 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1383 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1384 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1385 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1386 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1387 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1388 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1389 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1390 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1391 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1392 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1393 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1394 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1395 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1396 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1397 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1398 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1399 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1400 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1401 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1402 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1403 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1404 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1405 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1406 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1407 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1408 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1409 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1410 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1411 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1412 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1413 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1414 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1415 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1416 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1417 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1418 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1419 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1420 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1421 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1422 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1423 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1424 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1425 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1426 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1427 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1428 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1429 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1430 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1431 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1432 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1433 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1434 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1435 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1436 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1437 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1438 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1439 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1440 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1441 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1442 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1443 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1444 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1445 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1446 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1447 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1448 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1449 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1450 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1451 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1452 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1453 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1454 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1455 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1456 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1457 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1458 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1459 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1460 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1461 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1462 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1463 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1464 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1465 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1466 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1467 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1468 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1469 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1470 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1471 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1472 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1473 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1474 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1475 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1476 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1477 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1478 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1479 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1480 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1481 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1482 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1483 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1484 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1485 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1486 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1487 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1488 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1489 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1490 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1491 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1492 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1493 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1494 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1495 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1496 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1497 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1498 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1499 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1500 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1501 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1502 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1503 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1504 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1505 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1506 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1507 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1508 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1509 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1510 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1511 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1512 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1513 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1514 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1515 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1516 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1517 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1518 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1519 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1520 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1521 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1522 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1523 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1524 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1525 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1526 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1527 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1528 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1529 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1530 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1531 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1532 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1533 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1534 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1535 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1536 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1537 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1538 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1539 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1540 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1541 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1542 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1543 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1544 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1545 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1546 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1547 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1548 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1549 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1550 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1551 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1552 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1553 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1554 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1555 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1556 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1557 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1558 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1559 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1560 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1561 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1562 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1563 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1564 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1565 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1566 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1567 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1568 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1569 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1570 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1571 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1572 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1573 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1574 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1575 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1576 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1577 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1578 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1579 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1580 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1581 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1582 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1583 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1584 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1585 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1586 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1587 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1588 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1589 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1590 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1591 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1592 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1593 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1594 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1595 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1596 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1597 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1598 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1599 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1600 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1601 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1602 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1603 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1604 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1605 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1606 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1607 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1608 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1609 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1610 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1611 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1612 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1613 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1614 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1615 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1616 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1617 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1618 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1619 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1620 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1621 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1622 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1623 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1624 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1625 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1626 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1627 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1628 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1629 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1630 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1631 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1632 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1633 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1634 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1635 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1636 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1637 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1638 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1639 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1640 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1641 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1642 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1643 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1644 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1645 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1646 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1647 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1648 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1649 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1650 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1651 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1652 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1653 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1654 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1655 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1656 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1657 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1658 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1659 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1660 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1661 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1662 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1663 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1664 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1665 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1666 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1667 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1668 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1669 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1670 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1671 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1672 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1673 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1674 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1675 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1676 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1677 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1678 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1679 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1680 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1681 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1682 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1683 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1684 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1685 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1686 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1687 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1688 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1689 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1690 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1691 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1692 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1693 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1694 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1695 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1696 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1697 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1698 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1699 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1700 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1701 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1702 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1703 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1704 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1705 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1706 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1707 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1708 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1709 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1710 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1711 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1712 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1713 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1714 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1715 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1716 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1717 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1718 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1719 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1720 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1721 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1722 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1723 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1724 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1725 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1726 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1727 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1728 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1729 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1730 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1731 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1732 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1733 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1734 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1735 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1736 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1737 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1738 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1739 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1740 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1741 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1742 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1743 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1744 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1745 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1746 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1747 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1748 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1749 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1750 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1751 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1752 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1753 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1754 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1755 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1756 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1757 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1758 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1759 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1760 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1761 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1762 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1763 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1764 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1765 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1766 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1767 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1768 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1769 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1770 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1771 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1772 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1773 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1774 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1775 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1776 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1777 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1778 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1779 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1780 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1781 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1782 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1783 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1784 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1785 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1786 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1787 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1788 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1789 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1790 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1791 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1792 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1793 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1794 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1795 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1796 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1797 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1798 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1799 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1800 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1801 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1802 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1803 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1804 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1805 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1806 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1807 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1808 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1809 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1810 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1811 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1812 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1813 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1814 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1815 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1816 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1817 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1818 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1819 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1820 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1821 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1822 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1823 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1824 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1825 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1826 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1827 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1828 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1829 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1830 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1831 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1832 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1833 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1834 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1835 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1836 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1837 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1838 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1839 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1840 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1841 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1842 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1843 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1844 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1845 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1846 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1847 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1848 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1849 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1850 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1851 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1852 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1853 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1854 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1855 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1856 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1857 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1858 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1859 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1860 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1861 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1862 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1863 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1864 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1865 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1866 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1867 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1868 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1869 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1870 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1871 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1872 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1873 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1874 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1875 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1876 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1877 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1878 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1879 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1880 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1881 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1882 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1883 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1884 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1885 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1886 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1887 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1888 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1889 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1890 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1891 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1892 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1893 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1894 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1895 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1896 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1897 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1898 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1899 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1900 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1901 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1902 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1903 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1904 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1905 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1906 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1907 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1908 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1909 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1910 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1911 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1912 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1913 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1914 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1915 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1916 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1917 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1918 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1919 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1920 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1921 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1922 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1923 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1924 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1925 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1926 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1927 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1928 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1929 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1930 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1931 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1932 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1933 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1934 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1935 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1936 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1937 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1938 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1939 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1940 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1941 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1942 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1943 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1944 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1945 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1946 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1947 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1948 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1949 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1950 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1951 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1952 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1953 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1954 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1955 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1956 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1957 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1958 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1959 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1960 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1961 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1962 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1963 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1964 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1965 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1966 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1967 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1968 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1969 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1970 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1971 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1972 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1973 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1974 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1975 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1976 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1977 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1978 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1979 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1980 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1981 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1982 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1983 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1984 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1985 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1986 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1987 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1988 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1989 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1990 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1991 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1992 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1993 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1994 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1995 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1996 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1997 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1998 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  1999 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2000 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2001 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2002 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2003 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2004 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2005 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2006 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2007 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2008 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2009 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2010 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2011 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2012 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2013 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2014 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2015 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2016 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2017 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2018 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2019 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2020 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2021 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2022 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2023 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2024 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2025 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2026 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2027 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2028 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2029 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2030 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2031 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2032 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2033 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2034 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2035 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2036 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2037 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2038 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2039 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2040 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2041 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2042 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2043 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2044 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2045 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2046 ; write = 1; writedata [63:0]  = 64'h40092AF77DB8CC83; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        
        #10 address =  2047 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 
        
        #10 byteenable = 8'hF0; 
        #10 address =  2048 ; write = 1; writedata [63:0]  = 64'h4018F0329122D34E; byteenable = 8'h0F; 

        #10 byteenable = 8'hF0; 
	     
        #10 read = 1;

        #10000 $finish();
    end
endmodule

